module mc2 (
);
    
endmodule