// 
// {MODULE_NAME}_top.v 
//

module {MODULE_NAME}_top (
    // General Signals //
    // --------------- //
    input  logic                          clk                , // clock signal
    input  logic                          rst_n              , // active low reset

    // Input Controls // 
    // -------------- //

    // Input Data // 
    // ---------- //

    // Output Controls // 
    // --------------- // 

    // Output Data // 
    // ----------- //

);

// Local Parameters // 
// ---------------- //

// Internal Wires //
// -------------- //

// Internal Registers //
// ------------------ //

// Logic //
// ----- //

// FFs //
// --- //

endmodule

//|~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~|//
//|                                               |//
//| 1. Project  :  veri_env                       |//
//| 2. Author   :  Etay Sela                      |//
//| 3. Date     :  2025-01-09                     |//
//| 4. Version  :  v4.2.0                         |//
//|                                               |//
//|~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~|//
