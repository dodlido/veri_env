module gs (
);
    
endmodule