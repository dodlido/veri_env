module m1 (
   input wire clk,
   input wire rst_n
);















endmodule