module mc1 (
);
    
endmodule