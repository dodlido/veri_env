// 
// {MODULE_NAME}_top.v 
//

module {MODULE_NAME}_top (
    // General Signals //
    // --------------- //
    input  logic                          clk                , // clock signal
    input  logic                          rst_n              , // active low reset

    // Input Controls // 
    // -------------- //

    // Input Data // 
    // ---------- //

    // Output Controls // 
    // --------------- // 

    // Output Data // 
    // ----------- //

);

// Local Parameters // 
// ---------------- //

// Internal Wires //
// -------------- //

// Internal Registers //
// ------------------ //

// Logic //
// ----- //

// FFs //
// --- //

endmodule
